module fcu (
	ifc_fcu.dut d
	);

endmodule
