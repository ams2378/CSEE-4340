/**
* @filename  		counter.sv 
*
* @brief     		counter for credits avaible for neighboring router buffers
* @author   		ddl2126	<ddl2126@columbia.edu>
*	     		
*  	 
*/

module counter(
	ifc_counter.dut d
);

endmodule
