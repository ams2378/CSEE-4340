/**
* filename  		queue.sv 
* brief			Simple queue with width 5 and input data length of 16 bits     		
* authors   		Adil sadik <ams2378@columbia.edu>
* data creation		11/11/12	
* 
* 
*	 
*/


module queue (
	ifc_queue.dut d
);



endmodule
