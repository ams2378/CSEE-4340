/**
* @filename  		address_gen.sv 
*
* @brief     		Generates the direction to which data flits need to be sent, comparing current router address to destination address.

* @author   		Dechhin Lama	<ddl2126@columbia.edu>
*	     		
*  	 
*/

module address_gen (
		ifc_addr.dut d
		);

endmodule

