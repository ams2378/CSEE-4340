module xor_gate( a_i, b_i, out_o );

input a_i, b_i;
output out_o;

assign out_o = a_i ^ b_i; // bitwise xor

endmodule
