// adder
module adder (ifc.dut d);
 assign d.sum = d.a + d.b;
endmodule
