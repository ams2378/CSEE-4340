/**
* @filename  		count.sv 
*
* @brief     		counter for credits avaible for neighboring router buffers
* @author   		ddl2126	<ddl2126@columbia.edu>
*	     		
*  	 
*/

module counter(
	input incr_i,
	input decr_i, 

	output credit_en_o;	
)
