


module queue (

	input clk,
	input rst_n,
	input pop_req_i,
	input [15:0] data_i,		

	output [15:0] data_o
)
