/**
* filename  		fcu.sv 
* brief			Flow Control Unit- implements credit based flow control    		
* authors   		Adil sadik <ams2378@columbia.edu>
* data creation		11/11/12	
* 
* 
*	 
*/



module fcu (
	ifc_fcu.dut d
	);

endmodule
