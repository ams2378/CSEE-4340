/**
* @filename  		counter.sv 
*
* @brief     		Counter for credits avaible for neighboring router buffers
* @author   		Dechhin Lama	<ddl2126@columbia.edu>
*	     		
*  	 
*/

module counter(
	ifc_counter.dut d
);

endmodule
