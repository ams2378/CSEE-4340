/**
* @filename  		decoder_5_32.sv
*
* @brief     		decoder to decode read and write address
* @authors   		Dechhin Lama <ddl2126@columbia.edu>
*				 
*/

module decoder_5_32 ( decoder_i, decoder_o );

	input [4:0] decoder_i;
	output [31:0] decoder_o;

	logic [31:0] mid;
	
	always_comb begin
		case(decoder_i)
		
			5'd0:   mid = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
			5'd1:   mid = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
			5'd2:   mid = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
			5'd3:   mid = 32'b0000_0000_0000_0000_0000_0000_0000_1000;

			5'd4:   mid = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
			5'd5:   mid = 32'b0000_0000_0000_0000_0000_0000_0010_0000;
			5'd6:   mid = 32'b0000_0000_0000_0000_0000_0000_0100_0000;
			5'd7:   mid = 32'b0000_0000_0000_0000_0000_0000_1000_0000;
	
			5'd8:   mid = 32'b0000_0000_0000_0000_0000_0001_0000_0000;
			5'd9:   mid = 32'b0000_0000_0000_0000_0000_0010_0000_0000;
			5'd10:  mid = 32'b0000_0000_0000_0000_0000_0100_0000_0000;
			5'd11:  mid = 32'b0000_0000_0000_0000_0000_1000_0000_0000;

			5'd12:  mid = 32'b0000_0000_0000_0000_0001_0000_0000_0000;
			5'd13:  mid = 32'b0000_0000_0000_0000_0010_0000_0000_0000;
			5'd14:  mid = 32'b0000_0000_0000_0000_0100_0000_0000_0000;
			5'd15:  mid = 32'b0000_0000_0000_0000_1000_0000_0000_0000;

			5'd16:  mid = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
			5'd17:  mid = 32'b0000_0000_0000_0010_0000_0000_0000_0000;
			5'd18:  mid = 32'b0000_0000_0000_0100_0000_0000_0000_0000;
			5'd19:  mid = 32'b0000_0000_0000_1000_0000_0000_0000_0000;
			
			5'd20:  mid = 32'b0000_0000_0001_0000_0000_0000_0000_0000;
			5'd21:  mid = 32'b0000_0000_0010_0000_0000_0000_0000_0000;
			5'd22:  mid = 32'b0000_0000_0100_0000_0000_0000_0000_0000;
			5'd23:  mid = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
		
			5'd24:  mid = 32'b0000_0001_0000_0000_0000_0000_0000_0000;
			5'd25:  mid = 32'b0000_0010_0000_0000_0000_0000_0000_0000;
			5'd26:  mid = 32'b0000_0100_0000_0000_0000_0000_0000_0000;
			5'd27:  mid = 32'b0000_1000_0000_0000_0000_0000_0000_0000;
		
			5'd28:  mid = 32'b0001_0000_0000_0000_0000_0000_0000_0000;
			5'd29:  mid = 32'b0010_0000_0000_0000_0000_0000_0000_0000;
			5'd30:  mid = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
			5'd31:  mid = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
			default: mid = '0;
		endcase
	end
	
	assign decoder_o = mid;	

endmodule
