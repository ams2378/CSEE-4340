

module xbar (
	ifc_xbar.dut d
);

endmodule
