/*-----------------------------------------------------
Design Name : router
File Name   : router.sv
Function    : Top level file 

author	    : Dechhin Lama <ddl2126@columbia.edu>
*///-----------------------------------------------------


module router (
	ifc.dut d
	);

/*
 * instantiate the fcc */
/*fcc fcc_unit(
	
);*/

/*
 * instantiate the inputbuffers */
/*inputbuffer inputbuffer_unit(

);*/

/*
 * instantiate the arbiter */

/*
 * instantiate the fcu */

/*
 * instantiate the address generator */


/*
 * instantiate the xbar */

endmodule

