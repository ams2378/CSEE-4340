


module queue (
	ifc_queue.dut d
);



endmodule
