/**
* filename  		arbiter.sv 
* brief			Arbiter module for the router     		
* authors   		Adil sadik <ams2378@columbia.edu>
* date creation		11/11/12	
* 
* 
*	 
*/

module arbiter (
		ifc_arb.dut d
		);

endmodule


